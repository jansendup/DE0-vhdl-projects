library ieee;
use ieee.std_logic_1164.all;

entity uart is
	port(clk_i, reset_i : in std_logic);
end uart;